interface alu_if;
    logic [3:0] a, b;
    logic [1:0] op;
    logic [3:0] y;
    logic       carry;
endinterface
